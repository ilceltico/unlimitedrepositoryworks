library ieee;
use ieee.numeric_std.all;
use ieee.std_logic_1164.all;
use work.vga_package.all;

package HI_package is
	-- Constants declarations
	type spaceship_type is (ALIEN_1, ALIEN_2, ALIEN_3, RAND_ALIEN, PLAYER);
	
	-- Hitbox declaration
	type hitbox_type is record 
		up_left_x         : integer;
		up_left_y         : integer;
		size_x				: integer;
		size_y				: integer;
	end record;
	
	-- Spaceship declaration 	
	type spaceship is record
		ship_type      	: spaceship_type;
		hitbox				: hitbox_type;
		-- visible			: std_logic;
		exploding			: std_logic;
	end record;	

	type img_pixels_type is array(0 to 31, 0 to 31) of std_logic;
	
	type sprite_type is record 
		img_pixels				: img_pixels_type;
		color 					: color_type;
	end record;
	
	CONSTANT dummy_sprite: sprite_type := 
	(
		(
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000010000000000000000",
		"00000000000000001000000000000000",
		"00000000000000001000000000000000",
		"00000000000000001000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000"
		),
		COLOR_WHITE
	);
	
end package;