library ieee;
use ieee.numeric_std.all;
use ieee.std_logic_1164.all;
use work.vga_package.all;

package HI_package is

	-- Common constants
	constant REFERENCE_TIME_50MHz							: natural 	:= 50; -- Generates 1 microsecond, based on a 50MHz clock
	
	constant SPRITE_COUNT									: natural 	:= 26;
	constant ALIEN_SPRITE_COUNT							: natural	:= 3;
	constant BULLET_SPRITE_COUNT							: natural 	:= 4;
	constant SHIELD_SPRITE_COUNT							: natural 	:= 4;
	constant SPRITE_SIZE										: natural 	:= 32;
	constant MAX_HITBOX_SIZE								: natural 	:= 128;
	
	constant ALIENS_PER_COLUMN								: natural	:= 5;
	constant COLUMNS_PER_GRID 								: natural  	:= 11;
	constant SHIELD_COUNT									: natural  	:= 16;
	constant BULLET_COUNT									: natural 	:= 3;
	constant ALIEN_SIZE_X									: natural 	:= 26;
	constant ALIEN_SIZE_y									: natural 	:= 26;
	constant ALIEN_SPACING_X								: natural 	:= 8;
	constant ALIEN_SPACING_Y								: natural 	:= 15;
	constant SIDE_MARGIN 									: natural 	:= 10;
	constant TOP_MARGIN 										: natural 	:= 10;
	constant BOTTOM_MARGIN 									: natural	:= 10;
	constant RAND_ALIEN_SIZE_X 							: natural 	:= 46;
	constant RAND_ALIEN_SIZE_Y								: natural	:= 26;
	constant INDEX_1_MAX										: natural 	:= 16; 
	-- Set this last one to the maximum value between SHIELDS_COUNT, BULLET_COUNT and COLUMNS_PER_GRID
	
	constant FRAME_TIME_1us 								: natural := 16666; --60fps
	constant H_DISP											: natural := 640 - 128;
	constant V_DISP											: natural := 480;
	--constant EXPLOSION_TIME_50MHz 						: natural := 15000000;
	--constant RAND_ALIEN_EXPLOSION_TIME_50MHz 			: natural := 25000000;
	
	constant RAND_GEN_W										: natural := 16;
	
	-- Player
	constant PLAYER_MOVEMENT_TIME_1us					: natural := 16666; --30fps
	constant PLAYER_SIZE_X 									: natural := 30;
	constant PLAYER_SIZE_Y 									: natural := 18;
	constant PLAYER_START_X 								: natural := (H_DISP - PLAYER_SIZE_X) / 2;
	constant PLAYER_START_Y 								: natural := V_DISP - 4*PLAYER_SIZE_Y - BOTTOM_MARGIN;
	constant PLAYER_LIVES 									: natural := 3;
	constant PLAYER_SPEED 									: natural := 3;
	constant PLAYER_SPRITE_COUNT							: natural := 3;
	
	-- Bullets
	constant ALIEN_BULLET_SHAPE							: natural := 3; -- Number of alien bullets shapes
	constant ALIEN_BULLET_TIME_1us	 					: natural := 16666; --30 fps
	constant ALIEN_BULLET_SPEED 							: natural := 3;
	constant ALIEN_BULLET_SIZE_X 							: natural := 10;
	constant ALIEN_BULLET_SIZE_Y 							: natural := 20;
	constant PLAYER_BULLET_TIME_1us						: natural := 16666; --30 fps
	constant PLAYER_BULLET_SPEED 							: natural := 8;
	constant PLAYER_BULLET_SIZE_X 						: natural := 3;
	constant PLAYER_BULLET_SIZE_Y 						: natural := 8;
	constant BULLET_EXPLOSION_SIZE_X 					: natural := 30;
	constant BULLET_EXPLOSION_SIZE_Y 					: natural := 35;
	constant BULLET_EXPLOSION_TIME_50MHz 				: natural := 10000000;
	
	-- Alien points 
	constant ALIEN_1_POINTS 								: natural := 10;
	constant ALIEN_2_POINTS 								: natural := 20;
	constant ALIEN_3_POINTS 								: natural := 30;
	constant ALIEN_4_POINTS 								: natural := 300;
		
	-- Shields
	constant SHIELD_SIZE_X 									: natural := 33;
	constant SHIELD_SIZE_Y 									: natural := 33;
	constant SHIELD_SPACING 								: natural := 55;
	constant SHIELD_H_OVERLAP 								: natural := 7;
	constant SHIELD_V_OVERLAP 								: natural := 7;
	constant SHIELD_1_Y 										: natural := PLAYER_START_Y - SHIELD_SIZE_Y * 2 - 20;
	constant SHIELD_2_Y 										: natural := SHIELD_1_Y + SHIELD_SIZE_Y - SHIELD_V_OVERLAP;
	
	-- Level
	constant LEVEL_NUMBER 									: natural := 3;
	constant ALIEN_1_ROWS									: natural := 2;
	constant ALIEN_2_ROWS									: natural := 2;
	constant ALIEN_3_ROWS									: natural := 1;
	constant FIRST_ALIEN_CELL_X 							: natural := SIDE_MARGIN + 0;
	constant FIRST_ALIEN_CELL_Y 							: natural := TOP_MARGIN + RAND_ALIEN_SIZE_Y + 10;
	-- constant FIRST_RAND_ALIEN_CELL_X 					: natural := - RAND_ALIEN_SIZE_X;
	constant FIRST_RAND_ALIEN_CELL_X 					: integer := SIDE_MARGIN - RAND_ALIEN_SIZE_X;
	constant FIRST_RAND_ALIEN_CELL_Y 					: natural := TOP_MARGIN + 40;
	constant ALIEN_DOWN_SPEED 								: natural := 20;
	constant ALIEN_SPEED 									: natural := 10; --Aliens will be horizontally moved by this amount of pixels
	constant BASE_ALIEN_FRAME_TIME_1us	 				: natural := 1000000; --1fps
	constant ALIEN_FRAME_TIME_DECREASE_1us 			: natural := (BASE_ALIEN_FRAME_TIME_1us - FRAME_TIME_1us) / (ALIENS_PER_COLUMN * COLUMNS_PER_GRID - 1); -- Time decrease each time an alien gets destroyed
	constant BASE_ALIEN_BULLET_GEN_TIME_1us 		: natural := 2000000; --One bullet per 2 seconds
	--constant MAX_ALIEN_BULLET_GEN_TIME_50MHz 			: natural := 15000000; --More than 3 bullets per second
	--constant ALIEN_BULLET_GEN_TIME_DECREASE_50MHz 	: natural := (BASE_ALIEN_BULLET_GEN_TIME_50MHz - MAX_ALIEN_BULLET_GEN_TIME_50MHz) / (ALIENS_PER_COLUMN * COLUMNS_PER_GRID - 1);
	--constant BASE_ALIEN_BULLET_TIME_50MHz 				: natural := 50000000; --One bullet per second
	--constant MAX_ALIEN_BULLET_TIME_50MHz 				: natural := 15000000; --More than 3 bullets per second
	--constant ALIEN_BULLET_TIME_DECREASE_50MHz 		: natural := (BASE_ALIEN_BULLET_TIME_50MHz - MAX_ALIEN_BULLET_TIME_50MHz) / (ALIENS_PER_COLUMN * COLUMNS_PER_GRID - 1);
	constant RAND_ALIEN_SPEED 								: natural := 1;
	constant RAND_ALIEN_FRAME_TIME_1us 				: natural := 16666; --60fps
	constant RAND_ALIEN_TIME_RANGE_1us				: natural := 40000000; -- Time interval of 40 seconds
	constant RAND_ALIEN_TIME_MIN_1us					: natural := 20000000; -- Time interval of 20 seconds
	
	-- Sprites
	constant ALIEN_1_1_SPRITE 								: natural := 0;
	constant ALIEN_1_2_SPRITE 								: natural := 1;	 
	constant ALIEN_2_1_SPRITE 								: natural := 2;
	constant ALIEN_2_2_SPRITE 								: natural := 3;
	constant ALIEN_3_1_SPRITE 								: natural := 4;
	constant ALIEN_3_2_SPRITE 								: natural := 5;
	constant ALIEN_4_SPRITE  								: natural := 6;
	constant ALIEN_BULLET_1_1_SPRITE						: natural := 7;
	constant ALIEN_BULLET_1_2_SPRITE						: natural := 8;
	constant ALIEN_BULLET_1_3_SPRITE						: natural := 9;
	constant ALIEN_BULLET_1_4_SPRITE						: natural := 10;
	constant ALIEN_BULLET_2_1_SPRITE						: natural := 11;
	constant ALIEN_BULLET_2_2_SPRITE						: natural := 12;
	constant ALIEN_BULLET_2_3_SPRITE						: natural := 13;
	constant ALIEN_BULLET_2_4_SPRITE						: natural := 14;
	constant ALIEN_BULLET_3_1_SPRITE						: natural := 15;
	constant ALIEN_BULLET_3_2_SPRITE						: natural := 16;
	constant ALIEN_BULLET_3_3_SPRITE						: natural := 17;
	constant ALIEN_BULLET_3_4_SPRITE						: natural := 18;
	constant ALIEN_BULLET_EXPLOSION_SPRITE				: natural := 19;
	constant ALIEN_EXPLOSION_SPRITE						: natural := 20;
	constant PLAYER_SPRITE									: natural := 21;
	constant PLAYER_BULLET_SPRITE							: natural := 22;
	constant PLAYER_BULLET_EXPLOSION_SPRITE			: natural := 23;
	constant PLAYER_EXPLOSION_1_SPRITE					: natural := 24;
	constant PLAYER_EXPLOSION_2_SPRITE					: natural := 25;
	
	--------------------------------------------------------------
	--					            HITBOX				               --
	--------------------------------------------------------------
	
	-- Hitbox type declaration
	subtype hitbox_size is integer range 0 to MAX_HITBOX_SIZE - 1;
	type hitbox_type is record 
		up_left_x         : integer;
		up_left_y         : integer;
		size_x				: hitbox_size;
		size_y				: hitbox_size;
	end record;
	
	--------------------------------------------------------------
	--									SPRITE                           --
	--------------------------------------------------------------
	
	-- Sprite type declaration
	type img_pixels_type is array(0 to SPRITE_SIZE - 1 , 0 to SPRITE_SIZE - 1) of std_logic;
	subtype img_pixel_index_type is integer range 0 to SPRITE_SIZE - 1;
	subtype sprite_logic_dim_type is integer range 1 to SPRITE_SIZE;
	type sprite_type is record 
		img_pixels				: img_pixels_type;
		logic_dim_x				: sprite_logic_dim_type;
		logic_dim_y				: sprite_logic_dim_type;
		color 					: color_type;
	end record;
	
	-- Array of all sprites
	type sprite_array_type is array (0 to SPRITE_COUNT - 1) of sprite_type;
	subtype sprite_array_index_type is integer range 0 to SPRITE_COUNT - 1;
	
	constant sprite_empty : sprite_type := 
	(
		( 
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000"
		),
		32,
		32,
		COLOR_BLACK
	);
	
	--------------------------------------------------------------
	--	   							 PLAYER                          --
	--------------------------------------------------------------
	
	-- Player type declaration
	type player_sprite_indexes_type is array(0 to PLAYER_SPRITE_COUNT - 1) of sprite_array_index_type;
	subtype player_sprite_current_index_type is integer range 0 to PLAYER_SPRITE_COUNT - 1;
	subtype player_lives_type is integer range 0 to PLAYER_LIVES;
	type player_type is record
		sprite_indexes   	: player_sprite_indexes_type;
		hitbox				: hitbox_type;
		current_index		: player_sprite_current_index_type;
		lives					: player_lives_type;
		exploding			: std_logic;
	end record;	
	
	--------------------------------------------------------------
	--	   							 ALIEN                           --
	--------------------------------------------------------------
	
	-- Alien type declaration
	type alien_sprite_indexes_type is array(0 to ALIEN_SPRITE_COUNT - 1) of sprite_array_index_type;
	subtype alien_sprite_current_index_type is integer range 0 to ALIEN_SPRITE_COUNT - 1;
	type alien_type is record
		sprite_indexes   	: alien_sprite_indexes_type;
		hitbox				: hitbox_type;
		current_index		: alien_sprite_current_index_type;
		visible				: std_logic;
		exploding			: std_logic;
	end record;	
	
	-- Alien Column type declaration
	type alien_column_type is array(0 to ALIENS_PER_COLUMN - 1) of alien_type;
	subtype alien_column_index_type is integer range 0 to ALIENS_PER_COLUMN - 1;
	
	-- Alien Grid type declaration
	type alien_grid_type is array(0 to COLUMNS_PER_GRID - 1) of alien_column_type;
	subtype alien_grid_index_type is integer range 0 to COLUMNS_PER_GRID - 1;
	
	--------------------------------------------------------------
	--									BULLET                           --
	--------------------------------------------------------------
	
	-- Bullet type declaration
	type bullet_sprite_indexes_type is array(0 to BULLET_SPRITE_COUNT - 1) of sprite_array_index_type;
	subtype bullet_sprite_current_index_type is integer range 0 to BULLET_SPRITE_COUNT - 1;
	type bullet_type is record 
		sprite_indexes : bullet_sprite_indexes_type;
		hitbox			: hitbox_type;
		current_index	: bullet_sprite_current_index_type;
		visible			: std_logic;
		exploding		: std_logic;
	end record;
	
	-- Bullet array type declaration
	type bullet_array_type is array(0 to BULLET_COUNT - 1) of bullet_type;
	subtype bullet_array_index_type is integer range 0 to BULLET_COUNT - 1;
	
	subtype bullet_shape_type is integer range 0 to ALIEN_BULLET_SHAPE - 1;
	
	--------------------------------------------------------------
	--									SHIELD                           --
	--------------------------------------------------------------
	
	-- Shield type declaration
	type shield_sprite_indexes_type is array(0 to SHIELD_SPRITE_COUNT - 1) of sprite_array_index_type;
	subtype shield_sprite_current_index_type is integer range 0 to SHIELD_SPRITE_COUNT - 1;
	type shield_type is record 
		sprite_indexes : shield_sprite_indexes_type;
		hitbox			: hitbox_type;
		current_index	: shield_sprite_current_index_type;
		visible			: std_logic;
	end record;
	
	-- Bullet array type declaration
	type shield_array_type is array(0 to SHIELD_COUNT - 1) of shield_type;
	subtype shield_array_index_type is integer range 0 to SHIELD_COUNT - 1;
	
	--------------------------------------------------------------
	--					        DATAPATH INDEXES                     --
	--------------------------------------------------------------
	
	-- Datapath entity index type
	type entity_type_type is (ENTITY_NONE, ENTITY_ALIEN, ENTITY_ALIEN_BULLET, ENTITY_PLAYER_BULLET, ENTITY_SHIELD, ENTITY_RANDOM_ALIEN, ENTITY_PLAYER, ENTITY_COLUMN, ENTITY_BORDER);
	subtype index_1_type is integer range 0 to INDEX_1_MAX - 1;
	type datapath_entity_index_type is record
		index_1		: index_1_type;
		index_2 		: alien_column_index_type;
		entity_type : entity_type_type;
	end record;
	
	-- Datapath entity explosion index type
	type entity_explosion_index_type is record
		alien_row_index 			: alien_grid_index_type;
		alien_column_index 		: alien_column_index_type; 
		alien_exploding			: std_logic;
		
		bullet_index				: bullet_array_index_type;
		bullet_exploding			: std_logic;
		
		shield_index				: shield_array_index_type;
		shield_exploding			: std_logic;
		
		player_bullet_exploding : std_logic;
		player_exploding			: std_logic;
		random_alien_exploding	: std_logic;
	end record;
	
	type direction_type is (DIR_LEFT, DIR_RIGHT, DIR_UP, DIR_DOWN, DIR_NONE);
	
	--------------------------------------------------------------
	--					        DATAPATH INDEXES                     --
	--------------------------------------------------------------
	
	type collision_type is record 
		first_entity 			: datapath_entity_index_type;
		second_entity 			: datapath_entity_index_type;
	end record;
	
	--------------------------------------------------------------
	--					     ARRAY OF ALL SPRITES	                  --
	--------------------------------------------------------------	
	
-- 0 	-> Alien1_1.png
-- 1 	-> Alien1_2.png
-- 2 	-> Alien2_1.png
-- 3 	-> Alien2_2.png
-- 4 	-> Alien3_1.png
-- 5 	-> Alien3_2.png
-- 6 	-> Alien4.png
-- 7 	-> AlienBullet1_1.png
-- 8 	-> AlienBullet1_2.png
-- 9 	-> AlienBullet1_3.png
-- 10 -> AlienBullet1_4.png
-- 11 -> AlienBullet2_1.png
-- 12 -> AlienBullet2_2.png
-- 13 -> AlienBullet2_3.png
-- 14 -> AlienBullet2_4.png
-- 15 -> AlienBullet3_1.png
-- 16 -> AlienBullet3_2.png
-- 17 -> AlienBullet3_3.png
-- 18 -> AlienBullet3_4.png
-- 19 -> AlienBulletExplosion.png
-- 20 -> AlienExplosion.png
-- 21 -> Player.png
-- 22 -> PlayerBullet.png
-- 23 -> PlayerBulletExplosion.png
-- 24 -> PlayerExplosion1.png
-- 25 -> PlayerExplosion2.png
	
	constant sprites: sprite_array_type := 
	(
		-- 0 	-> Alien1_1.png
		(
			( 
				"00001111000000000000000000000000",
				"01111111111000000000000000000000",
				"11111111111100000000000000000000",
				"11100110011100000000000000000000",
				"11111111111100000000000000000000",
				"00011001100000000000000000000000",
				"00100110010000000000000000000000",
				"00010000100000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000"
			),
			12,
			8,
			COLOR_WHITE
		),
		-- 1 	-> Alien1_2.png
		(	
			( 
				"00001111000000000000000000000000",
				"01111111111000000000000000000000",
				"11111111111100000000000000000000",
				"11100110011100000000000000000000",
				"11111111111100000000000000000000",
				"00011001100000000000000000000000",
				"00110110110000000000000000000000",
				"11000000001100000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000"
			),
			12,
			8,
			COLOR_WHITE
		),
		-- 2 	-> Alien2_1.png
		( 
			(
				"00100000100000000000000000000000",
				"00010001000000000000000000000000",
				"00111111100000000000000000000000",
				"01101110110000000000000000000000",
				"11111111111000000000000000000000",
				"10111111101000000000000000000000",
				"10100000101000000000000000000000",
				"00011011000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000"
			),
			11,
			8,
			COLOR_WHITE
		),
		-- 3 	-> Alien2_2.png
		( 
			(
				"00100000100000000000000000000000",
				"10010001001000000000000000000000",
				"10111111101000000000000000000000",
				"11101110111000000000000000000000",
				"11111111111000000000000000000000",
				"00111111100000000000000000000000",
				"00100000100000000000000000000000",
				"01000000010000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000"
			),
			11,
			8,
			COLOR_WHITE
		),
		-- 4 	-> Alien3_1.png
		( 
			(
				"00011000000000000000000000000000",
				"00111100000000000000000000000000",
				"01111110000000000000000000000000",
				"11011011000000000000000000000000",
				"11111111000000000000000000000000",
				"00100100000000000000000000000000",
				"01011010000000000000000000000000",
				"10100101000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000"
			),
			8,
			8,
			COLOR_WHITE
		),
		-- 5 	-> Alien3_2.png
		( 
			(
				"00011000000000000000000000000000",
				"00111100000000000000000000000000",
				"01111110000000000000000000000000",
				"11011011000000000000000000000000",
				"11111111000000000000000000000000",
				"00100100000000000000000000000000",
				"01000010000000000000000000000000",
				"00100100000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000"
			),
			8,
			8,
			COLOR_WHITE
		),
		-- 6 	-> Alien4.png
		( 
			(
				"00000111111000000000000000000000",
				"00011111111110000000000000000000",
				"00111111111111000000000000000000",
				"01101101101101100000000000000000",
				"11111111111111110000000000000000",
				"00111001100111000000000000000000",
				"00010000000010000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000"
			),
			16,
			7,
			COLOR_WHITE
		),
		-- 7 	-> AlienBullet1_1.png
		( 
			(
				"10000000000000000000000000000000",
				"10000000000000000000000000000000",
				"10000000000000000000000000000000",
				"10000000000000000000000000000000",
				"10000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000"
			),
			1,
			5,
			COLOR_WHITE
		),
		-- 8 	-> AlienBullet1_2.png
		( 
			(
				"01111000000000000000000000000000",
				"11111000000000000000000000000000",
				"11110000000000000000000000000000",
				"11110000000000000000000000000000",
				"01111000000000000000000000000000",
				"01111000000000000000000000000000",
				"11111000000000000000000000000000",
				"11111000000000000000000000000000",
				"11110000000000000000000000000000",
				"01110000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000"
			),
			5,
			10,
			COLOR_WHITE
		),
		-- 9 	-> AlienBullet1_3.png
		( 
			(
				"01110000000000000000000000000000",
				"01110000000000000000000000000000",
				"01110000000000000000000000000000",
				"01110000000000000000000000000000",
				"01110000000000000000000000000000",
				"01110000000000000000000000000000",
				"01110000000000000000000000000000",
				"01110000000000000000000000000000",
				"01110000000000000000000000000000",
				"01110000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000"
			),
			4,
			10,
			COLOR_WHITE
		),
		-- 10 -> AlienBullet1_4.png
		( 
			(
				"01110000000000000000000000000000",
				"01111000000000000000000000000000",
				"11111000000000000000000000000000",
				"11111000000000000000000000000000",
				"11110000000000000000000000000000",
				"11110000000000000000000000000000",
				"01111000000000000000000000000000",
				"01111000000000000000000000000000",
				"11111000000000000000000000000000",
				"11110000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000"
			),
			5,
			10,
			COLOR_WHITE
		),
		-- 11 -> AlienBullet2_1.png
		( 
			(
				"11110000000000000000000000000000",
				"11111100000000000000000000000000",
				"01111100000000000000000000000000",
				"01111100000000000000000000000000",
				"11111000000000000000000000000000",
				"11111000000000000000000000000000",
				"01111100000000000000000000000000",
				"01111100000000000000000000000000",
				"01111100000000000000000000000000",
				"11111000000000000000000000000000",
				"11110000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000"
			),
			6,
			11,
			COLOR_WHITE
		),
		-- 12 -> AlienBullet2_2.png
		( 
			(
				"00111100000000000000000000000000",
				"11111100000000000000000000000000",
				"11111000000000000000000000000000",
				"11111000000000000000000000000000",
				"01111100000000000000000000000000",
				"01111100000000000000000000000000",
				"11111000000000000000000000000000",
				"11111000000000000000000000000000",
				"11111000000000000000000000000000",
				"01111100000000000000000000000000",
				"00111100000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000"
			),
			6,
			11,
			COLOR_WHITE
		),
		-- 13 -> AlienBullet2_3.png
		( 
			(
				"11100000000000000000000000000000",
				"11111000000000000000000000000000",
				"01111100000000000000000000000000",
				"01111100000000000000000000000000",
				"01111100000000000000000000000000",
				"01111000000000000000000000000000",
				"11111000000000000000000000000000",
				"11110000000000000000000000000000",
				"01110000000000000000000000000000",
				"01111100000000000000000000000000",
				"00011100000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000"
			),
			6,
			11,
			COLOR_WHITE
		),
		-- 14 -> AlienBullet2_4.png
		( 
			(
				"11110000000000000000000000000000",
				"11111100000000000000000000000000",
				"01111100000000000000000000000000",
				"01111100000000000000000000000000",
				"11111000000000000000000000000000",
				"11111000000000000000000000000000",
				"01111100000000000000000000000000",
				"01111100000000000000000000000000",
				"01111100000000000000000000000000",
				"11111000000000000000000000000000",
				"11110000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000"
			),
			6,
			11,
			COLOR_WHITE
		),
		-- 15 -> AlienBullet3_1.png
		( 
			(
				"11111000000000000000000000000000",
				"11111000000000000000000000000000",
				"01110000000000000000000000000000",
				"01110000000000000000000000000000",
				"01110000000000000000000000000000",
				"01110000000000000000000000000000",
				"01110000000000000000000000000000",
				"01110000000000000000000000000000",
				"01110000000000000000000000000000",
				"01110000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000"
			),
			5,
			10,
			COLOR_WHITE
		),
		-- 16 -> AlienBullet3_2.png
		( 
			(
				"01110000000000000000000000000000",
				"11111000000000000000000000000000",
				"11111000000000000000000000000000",
				"11111000000000000000000000000000",
				"01110000000000000000000000000000",
				"01110000000000000000000000000000",
				"01110000000000000000000000000000",
				"01110000000000000000000000000000",
				"01110000000000000000000000000000",
				"01110000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000"
			),
			5,
			10,
			COLOR_WHITE
		),
		-- 17 -> AlienBullet3_3.png
		( 
			(
				"01110000000000000000000000000000",
				"01110000000000000000000000000000",
				"01110000000000000000000000000000",
				"01110000000000000000000000000000",
				"01110000000000000000000000000000",
				"11111000000000000000000000000000",
				"11111000000000000000000000000000",
				"11111000000000000000000000000000",
				"01110000000000000000000000000000",
				"01110000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000"
			),
			5,
			10,
			COLOR_WHITE
		),
		-- 18 -> AlienBullet3_4.png
		( 
			(
				"01110000000000000000000000000000",
				"01110000000000000000000000000000",
				"01110000000000000000000000000000",
				"01110000000000000000000000000000",
				"01110000000000000000000000000000",
				"01110000000000000000000000000000",
				"01110000000000000000000000000000",
				"01110000000000000000000000000000",
				"11111000000000000000000000000000",
				"11111000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000"
			),
			5,
			10,
			COLOR_WHITE
		),
		-- 19 -> AlienBulletExplosion.png
		( 
			(
				"00000000000000111000000000000000",
				"00000000000000111000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000001110000000000",
				"00000000001110000001110000000000",
				"00000000001110000001100000000000",
				"00000000001111110000000000000000",
				"00000011100001111110000000111000",
				"00000011100001111110000000111000",
				"00000011100001111100111000111000",
				"00000000001101111111111110000000",
				"00000000001111111111111110000000",
				"00000000001111111111111110000000",
				"00000001111111111111111111100000",
				"00011101111111101111111111100000",
				"00011011111111111111111111111100",
				"00011111111111111111111111111100",
				"00001110011111111111111111000000",
				"00001110001111111111111111000000",
				"11000000000011111111111111000000",
				"11000000001111110011011111000000",
				"11000000001110111111011000000000",
				"00000000000000001111100001110000",
				"00000000000000000001100001110000",
				"00000000001110000001100001100000",
				"00000000001110000000000000000000",
				"00000000000001100000000000000000",
				"00000000000001100000000000000000",
				"00000000000001100000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000"
			),
			32,
			29,
			COLOR_WHITE
		),
		-- 20 -> AlienExplosion.png
		( 
			(
				"00000011000001100000000000000000",
				"01100011000001100011000000000000",
				"01100000110110000011000000000000",
				"00011000110110001100000000000000",
				"00011110000000111100000000000000",
				"00000110000000110000000000000000",
				"11110000000000000111100000000000",
				"11110110000000110111100000000000",
				"00000110000000110000000000000000",
				"00011000110110001100000000000000",
				"00011011110111101100000000000000",
				"01100011000001100111000000000000",
				"01100000000000000010000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000"
			),
			21,
			13,
			COLOR_WHITE
		),
		-- 21 -> Player.png
		( 
			(
				"00000010000000000000000000000000",
				"00000111000000000000000000000000",
				"00000111000000000000000000000000",
				"01111111111100000000000000000000",
				"11111111111110000000000000000000",
				"11111111111110000000000000000000",
				"11111111111110000000000000000000",
				"11111111111110000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000"
			),
			13,
			8,
			COLOR_WHITE
		),
		-- 22 -> PlayerBullet.png
		( 
			(
				"11000000000000000000000000000000",
				"11000000000000000000000000000000",
				"11000000000000000000000000000000",
				"11000000000000000000000000000000",
				"11000000000000000000000000000000",
				"11000000000000000000000000000000",
				"11000000000000000000000000000000",
				"11000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000"
			),
			2,
			8,
			COLOR_WHITE
		),
		-- 23 -> PlayerBulletExplosion.png
		( 
			(
				"00000000001110000000000000000000",
				"00000000011110000000000000000000",
				"00000000011110000001110000000000",
				"00000000011110011001110000000000",
				"00000000001001111001110000000000",
				"00111000001101111000000000000000",
				"00111000111111111110000111000000",
				"00111000111111111110011110000000",
				"00000000111111111111111111100000",
				"00000111111111111111111111100000",
				"00000111111111111111100011100000",
				"00111111111111111111110000000000",
				"11111001111111111111110000000000",
				"11111000011111111111110000000000",
				"11100000011111111111100000000000",
				"00000000011111111111100000000000",
				"00000011111111111111001110000000",
				"00000111111011111110001110000000",
				"00000111111000111000001110000000",
				"00000000001110000000000000000000",
				"00000000001110001100000000000000",
				"00000000001110001110000000000000",
				"00000000000000001110000000000000",
				"00000000000000001100000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000"
			),
			27,
			24,
			COLOR_WHITE
		),
		-- 24 -> PlayerExplosion1.png
		( 
			(
				"00000100000000000000000000000000",
				"00000000001000000000000000000000",
				"00000101010000000000000000000000",
				"00100100000000000000000000000000",
				"00000011011000000000000000000000",
				"10001011010100000000000000000000",
				"00111111110010000000000000000000",
				"01111111111010100000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000"
			),
			15,
			8,
			COLOR_WHITE
		),
		-- 25 -> PlayerExplosion2.png
		( 
			(
				"00010000000001000000000000000000",
				"10000010000110010000000000000000",
				"00010000110000000000000000000000",
				"00000010000000100000000000000000",
				"01001011001100010000000000000000",
				"00100001110001000000000000000000",
				"00011111111100000000000000000000",
				"00110111111100100000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000",
				"00000000000000000000000000000000"
			),
			16,
			8,
			COLOR_WHITE
		)
	);
end package;