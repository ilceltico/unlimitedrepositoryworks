library ieee;
use ieee.numeric_std.all;
use ieee.std_logic_1164.all;
use work.vga_package.all;

package HI_package is
	-- Constants declarations
	constant ALIEN_SPRITE_COUNT	: positive	:= 3;
	constant ALIENS_PER_COLUMN		: positive	:= 1;
	constant COLUMNS_PER_GRID 		: positive  := 2;
	constant SPRITE_SIZE				: positive 	:= 32;
	
	
	-- Hitbox declaration
	type hitbox_type is record 
		up_left_x         : integer;
		up_left_y         : integer;
		size_x				: integer;
		size_y				: integer;
	end record;
	
	-- Spaceship declaration 	
	type alien_sprite_indexes_type is array(0 to ALIEN_SPRITE_COUNT - 1) of integer;
	subtype alien_sprite_current_index_type is integer range 0 to ALIEN_SPRITE_COUNT - 1;
	type alien_type is record
		sprite_indexes   	: alien_sprite_indexes_type;
		hitbox				: hitbox_type;
		current_index		: alien_sprite_current_index_type;
		-- visible			: std_logic;
		-- exploding		: std_logic;
	end record;	
	
	-- Alien Column declaration
	type alien_column_type is array(0 to ALIENS_PER_COLUMN - 1) of alien_type;
	subtype alien_column_index_type is integer range 0 to ALIENS_PER_COLUMN - 1;
	
	-- Alien Grid declaration
	type alien_grid_type is array(0 to COLUMNS_PER_GRID - 1) of alien_column_type;
	subtype alien_grid_index_type is integer range 0 to COLUMNS_PER_GRID - 1;
	

	type img_pixels_type is array(0 to SPRITE_SIZE - 1 , 0 to SPRITE_SIZE - 1) of std_logic;
	subtype img_pixel_index_type is integer range 0 to SPRITE_SIZE - 1;
	
	type sprite_type is record 
		img_pixels				: img_pixels_type;
		logic_dim_x				: integer;
		logic_dim_y				: integer;
		color 					: color_type;
	end record;
	
	type sprite_array_type is array (0 to 2) of sprite_type;
	
	constant sprites: sprite_array_type := 
	(
		(
			(
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000011100000000000000111000000",
			"00000011100000000000000111000000",
			"00000011100000000000000111000000",
			"00000000011100000000111000000000",
			"00000000011100000000111000000000",
			"00000000011100000000111000000000",
			"00000011111111111111111111000000",
			"00000011111111111111111111000000",
			"00000011111111111111111111000000",
			"00011111100011111111000111111000",
			"00011111100011111111000111111000",
			"00011111100011111111000111111000",
			"11111111111111111111111111111111",
			"11111111111111111111111111111111",
			"11111111111111111111111111111111",
			"11100011111111111111111111000111",
			"11100011111111111111111111000111",
			"11100011111111111111111111000111",
			"11100011100000000000000111000111",
			"11100011100000000000000111000111",
			"11100011100000000000000111000111",
			"00000000011111100111111000000000",
			"00000000011111100111111000000000",
			"00000000011111100111111000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000"
			),
			32,
			32,
			COLOR_WHITE
		),
		(	
			(
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000011100000000000000111000000",
			"00000011100000000000000111000000",
			"00000011100000000000000111000000",
			"11100000011100000000111000000111",
			"11100000011100000000111000000111",
			"11100000011100000000111000000111",
			"11100011111111111111111111000111",
			"11100011111111111111111111000111",
			"11100011111111111111111111000111",
			"11111111100011111111000111111111",
			"11111111100011111111000111111111",
			"11111111100011111111000111111111",
			"11111111111111111111111111111111",
			"11111111111111111111111111111111",
			"11111111111111111111111111111111",
			"00011111111111111111111111111000",
			"00011111111111111111111111111000",
			"00011111111111111111111111111000",
			"00000011100000000000000111000000",
			"00000011100000000000000111000000",
			"00000011100000000000000111000000",
			"00011100000000000000000000111000",
			"00011100000000000000000000111000",
			"00011100000000000000000000111000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000"
			),
			32,
			32,
			COLOR_WHITE
		),
		( 
			(
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000001110000001110000000000",
			"00011100011110000001110000111000",
			"00011100001111100111110000111000",
			"00011100000011100111000000111000",
			"00000111100011100111000111000000",
			"00000111100000000000000111000000",
			"00000000111000000000011100000000",
			"00000000111000000000011100000000",
			"00111110111000000000011101111100",
			"00111110000000000000000001111100",
			"00111110111000000000011101111100",
			"00000000111000000000011100000000",
			"00000000111011100111011100000000",
			"00000011100011100111000111000000",
			"00000011101111100111110111000000",
			"00011100011110000001110000111000",
			"00011100011110000001110000111000",
			"00011100000000000000000000111000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000"
			),
			32,
			32,
			COLOR_WHITE
		)
	);
end package;