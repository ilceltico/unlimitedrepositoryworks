library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity SpaceInvadersUnlimited is
		Port 
		( 
				CLOCK : in  std_logic;
				RESET : in  std_logic
		);
end entity;

architecture RTL of SpaceInvadersUnlimited is
	signal clock              : std_logic;

begin
end architecture;