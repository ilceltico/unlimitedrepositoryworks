library ieee;
use ieee.numeric_std.all;
use ieee.std_logic_1164.all;
use work.vga_package.all;

package HI_package is
	-- Constants declarations
	
	
	
	-- Hitbox declaration
	type hitbox_type is record 
		up_left_x         : integer;
		up_left_y         : integer;
		size_x				: integer;
		size_y				: integer;
	end record;
	
	-- Spaceship declaration 	
	type alien_sprite_indexes_type is array(0 to 2) of integer;
	subtype alien_sprite_current_index_type is integer range 0 to 2;
	type alien_type is record
		sprite_indexes   	: alien_sprite_indexes_type;
		hitbox				: hitbox_type;
		current_index		: alien_sprite_current_index_type;
		-- visible			: std_logic;
		-- exploding		: std_logic;
	end record;	

	type img_pixels_type is array(0 to 31, 0 to 31) of std_logic;
	
	
	type sprite_type is record 
		img_pixels				: img_pixels_type;
		color 					: color_type;
	end record;
	
	type sprite_array_type is array (0 to 1) of sprite_type;
	
	CONSTANT sprites: sprite_array_type := 
	(
		(
			(
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000111000000000001110000000",
			"00000000111000000000001110000000",
			"00000000000110000000110000000000",
			"00000000000110000000110000000000",
			"00000000011111111111111100000000",
			"00000000111111111111111110000000",
			"00000000111111111111111110000000",
			"00000011111001111111001111100000",
			"00000011111001111111001111100000",
			"00001111111111111111111111110000",
			"00001111111111111111111111110000",
			"00001100111111111111111110010000",
			"00001100111111111111111110010000",
			"00001100111111111111111110010000",
			"00001100111000000000001110010000",
			"00001100011000000000001100010000",
			"00000000000111110111110000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000"
			),
			COLOR_WHITE
		),
		(	
			(
			"11111111111111111111111111111111",
			"11111111111111111111111111111111",
			"11111111111111111111111111111111",
			"11111111110000000000000011111111",
			"11111111111111111111111111111111",
			"11111111111111111111111111111111",
			"11111111111111111111111111111111",
			"11111111111111111111111111111111",
			"11111111111111111111111111111111",
			"11111111111111111111111111111111",
			"11111111111111111111111111111111",
			"11111111111111111111111111111111",
			"11111111111111111111111111111111",
			"11111111111111111111111111111111",
			"11111111111111111111111111111111",
			"11111111111111111111111111111111",
			"11111111111111111111111111111111",
			"11111111111111111111111111111111",
			"11111111111111111111111111111111",
			"11111111111111111111111111111111",
			"11111111111111111111111111111111",
			"11111111111111111111111111111111",
			"11111111111111111111111111111111",
			"11111111111111111111111111111111",
			"11111111111111111111111111111111",
			"11111111111111111111111111111111",
			"11111111111111111111111111111111",
			"11111111111111111111111111111111",
			"11111111111111111111111111111111",
			"11111111111111111111111111111111",
			"11111111111111111111111111111111",
			"11111111111111111111111111111111"
			),
			COLOR_RED
		)
	);
end package;