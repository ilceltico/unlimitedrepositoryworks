-- source: https://www.nandland.com/vhdl/modules/double-dabble.html
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
 
entity Binary_to_BCD is
	generic (
		g_INPUT_WIDTH    : in positive := 15;
		g_DECIMAL_DIGITS : in positive := 4
   );
	port (
		CLOCK  : in std_logic;
		START  : in std_logic;
		BINARY : in std_logic_vector(g_INPUT_WIDTH-1 downto 0);
     
		o_BCD : out std_logic_vector(g_DECIMAL_DIGITS*4-1 downto 0);
		o_DV  : out std_logic
   );
end entity Binary_to_BCD;
 
architecture rtl of Binary_to_BCD is
 
	type t_BCD_State is (s_IDLE, s_SHIFT, s_CHECK_SHIFT_INDEX, s_ADD, s_CHECK_DIGIT_INDEX, s_BCD_DONE);
	signal r_SM_Main : t_BCD_State := s_IDLE;
 
	-- The vector that contains the output BCD
	signal r_BCD : std_logic_vector(g_DECIMAL_DIGITS*4-1 downto 0) := (others => '0');
 
	-- The vector that contains the input binary value being shifted.
	signal r_Binary : std_logic_vector(g_INPUT_WIDTH-1 downto 0) := (others => '0');
   
	-- Keeps track of which Decimal Digit we are indexing
	signal r_Digit_Index : natural range 0 to g_DECIMAL_DIGITS-1 := 0;
 
	-- Keeps track of which loop iteration we are on.
	-- Number of loops performed = g_INPUT_WIDTH
	signal r_Loop_Count : natural range 0 to g_INPUT_WIDTH-1  := 0;
   
begin
 
	Double_Dabble : process (CLOCK)
		variable v_Upper     : natural;
		variable v_Lower     : natural;
		variable mask			: std_logic_vector(g_DECIMAL_DIGITS*4-1 downto 0);
		variable r_BCD_temp	: std_logic_vector(g_DECIMAL_DIGITS*4-1 downto 0);
		variable v_BCD_Digit : unsigned(3 downto 0);
	begin
		if rising_edge(CLOCK) then
 
			case r_SM_Main is
 
			-- Stay in this state until i_Start comes along
			when s_IDLE =>
				if START = '1' then
					r_BCD     <= (others => '0');
					r_Binary  <= BINARY;
					r_SM_Main <= s_SHIFT;
				else
					r_SM_Main <= s_IDLE;
				end if;
 
			-- Always shift the BCD Vector until we have shifted all bits through
			-- Shift the most significant bit of r_Binary into r_BCD lowest bit.
			when s_SHIFT =>
				r_BCD     <= r_BCD(r_BCD'left-1 downto 0) & r_Binary(r_Binary'left);
				r_Binary  <= r_Binary(r_Binary'left-1 downto 0) & '0';
				r_SM_Main <= s_CHECK_SHIFT_INDEX;
 
			-- Check if we are done with shifting in r_Binary vector
			when s_CHECK_SHIFT_INDEX => 
				if r_Loop_Count = g_INPUT_WIDTH-1 then
					r_Loop_Count <= 0;
					r_SM_Main    <= s_BCD_DONE;
				else
					r_Loop_Count <= r_Loop_Count + 1;
					r_SM_Main    <= s_ADD;
				end if;
 
			-- Break down each BCD Digit individually.  Check them one-by-one to
			-- see if they are greater than 4. If they are, increment by 3.
			-- Put the result back into r_BCD Vector.  Note that v_BCD_Digit is
			-- unsigned.  Numeric_std does not perform math on std_logic_vector.
			when s_ADD =>
				
				v_Lower     := r_Digit_Index*4;
			
				mask 			:= (others => '0');
				mask(3 downto 0) := "1111";
				mask 			:= std_logic_vector(shift_left(unsigned(mask), v_Lower));
				mask 			:= mask and r_BCD;
				mask 			:= std_logic_vector(shift_right(unsigned(mask), v_Lower));
				
				v_BCD_Digit := unsigned(mask(3 downto 0));
           
				if v_BCD_Digit > 4 then
					v_BCD_Digit := v_BCD_Digit + 3;
				end if;
	
				mask 			:= (others => '0');
				mask(3 downto 0) := "1111";
				mask 			:= std_logic_vector(shift_left(unsigned(mask), v_Lower));
				mask 			:= not(mask);
				r_BCD_temp 	:= r_BCD;
				r_BCD_temp	:= r_BCD_temp and mask;
				mask 			:= (others => '0');
				mask(3 downto 0) := std_logic_vector(v_BCD_Digit);
				mask 			:= std_logic_vector(shift_left(unsigned(mask), v_Lower));
				r_BCD_temp	:= r_BCD_temp or mask;
				
				r_BCD <= r_BCD_temp;
		
				r_SM_Main <= s_CHECK_DIGIT_INDEX;
 
			-- Check if we are done incrementing all of the BCD Digits
			when s_CHECK_DIGIT_INDEX =>
				if r_Digit_Index = g_DECIMAL_DIGITS-1 then
					r_Digit_Index <= 0;
					r_SM_Main     <= s_SHIFT;
				else
					r_Digit_Index <= r_Digit_Index + 1;
					r_SM_Main     <= s_ADD;
				end if;
 
			when s_BCD_DONE =>
				r_SM_Main <= s_IDLE;
       
			when others =>
				r_SM_Main <= s_IDLE;
           
			end case;
		end if;            
	end process Double_Dabble;
 
	o_DV  <= '1' when r_SM_Main = s_BCD_DONE else '0';
	o_BCD <= r_BCD;
   
end architecture rtl;