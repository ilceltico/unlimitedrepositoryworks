library ieee;
  use ieee.std_logic_1164.all;
	use ieee.numeric_std.ALL;
    
package rand_gen_package is
    constant rand_gen_w : natural := 4;		-- LFSR width
end;