-- qsys.vhd

-- Generated using ACDS version 13.0sp1 232 at 2018.09.12.19:59:53

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity qsys is
	port (
		onchip_memory2_0_s1_address       : in  std_logic_vector(12 downto 0) := (others => '0'); --     onchip_memory2_0_s1.address
		onchip_memory2_0_s1_debugaccess   : in  std_logic                     := '0';             --                        .debugaccess
		onchip_memory2_0_s1_clken         : in  std_logic                     := '0';             --                        .clken
		onchip_memory2_0_s1_chipselect    : in  std_logic                     := '0';             --                        .chipselect
		onchip_memory2_0_s1_write         : in  std_logic                     := '0';             --                        .write
		onchip_memory2_0_s1_readdata      : out std_logic_vector(15 downto 0);                    --                        .readdata
		onchip_memory2_0_s1_writedata     : in  std_logic_vector(15 downto 0) := (others => '0'); --                        .writedata
		onchip_memory2_0_s1_byteenable    : in  std_logic_vector(1 downto 0)  := (others => '0'); --                        .byteenable
		onchip_memory2_0_reset1_reset     : in  std_logic                     := '0';             -- onchip_memory2_0_reset1.reset
		onchip_memory2_0_reset1_reset_req : in  std_logic                     := '0';             --                        .reset_req
		onchip_memory2_0_clk1_clk         : in  std_logic                     := '0'              --   onchip_memory2_0_clk1.clk
	);
end entity qsys;

architecture rtl of qsys is
	component qsys_onchip_memory2_0 is
		port (
			clk         : in  std_logic                     := 'X';             -- clk
			address     : in  std_logic_vector(12 downto 0) := (others => 'X'); -- address
			debugaccess : in  std_logic                     := 'X';             -- debugaccess
			clken       : in  std_logic                     := 'X';             -- clken
			chipselect  : in  std_logic                     := 'X';             -- chipselect
			write       : in  std_logic                     := 'X';             -- write
			readdata    : out std_logic_vector(15 downto 0);                    -- readdata
			writedata   : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			byteenable  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable
			reset       : in  std_logic                     := 'X';             -- reset
			reset_req   : in  std_logic                     := 'X'              -- reset_req
		);
	end component qsys_onchip_memory2_0;

begin

	onchip_memory2_0 : component qsys_onchip_memory2_0
		port map (
			clk         => onchip_memory2_0_clk1_clk,         --   clk1.clk
			address     => onchip_memory2_0_s1_address,       --     s1.address
			debugaccess => onchip_memory2_0_s1_debugaccess,   --       .debugaccess
			clken       => onchip_memory2_0_s1_clken,         --       .clken
			chipselect  => onchip_memory2_0_s1_chipselect,    --       .chipselect
			write       => onchip_memory2_0_s1_write,         --       .write
			readdata    => onchip_memory2_0_s1_readdata,      --       .readdata
			writedata   => onchip_memory2_0_s1_writedata,     --       .writedata
			byteenable  => onchip_memory2_0_s1_byteenable,    --       .byteenable
			reset       => onchip_memory2_0_reset1_reset,     -- reset1.reset
			reset_req   => onchip_memory2_0_reset1_reset_req  --       .reset_req
		);

end architecture rtl; -- of qsys
